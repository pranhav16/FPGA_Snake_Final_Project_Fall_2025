library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity poison_control is
    generic (
        GRID_WIDTH    : integer := 40;
        GRID_HEIGHT   : integer := 30;
        VISIBLE_TICKS : integer := 80;
        HIDDEN_TICKS  : integer := 30;
        SEED          : std_logic_vector(9 downto 0) := "1100110011"
    );
    port (
        clk       : in  std_logic;
        rst       : in  std_logic;
        game_tick : in  std_logic;
        p1_head_x : in  integer range 0 to GRID_WIDTH-1;
        p1_head_y : in  integer range 0 to GRID_HEIGHT-1;
        p2_head_x : in  integer range 0 to GRID_WIDTH-1;
        p2_head_y : in  integer range 0 to GRID_HEIGHT-1;

        -- dynamic walls (from wall_field)
        w1_x0_i        : in integer range 0 to GRID_WIDTH-1;
        w1_y0_i        : in integer range 0 to GRID_HEIGHT-1;
        w1_orient_i    : in std_logic;
        w2_x0_i        : in integer range 0 to GRID_WIDTH-1;
        w2_y0_i        : in integer range 0 to GRID_HEIGHT-1;
        w2_orient_i    : in std_logic;
        w3_x0_i        : in integer range 0 to GRID_WIDTH-1;
        w3_y0_i        : in integer range 0 to GRID_HEIGHT-1;
        w3_orient_i    : in std_logic;
        walls_solid_i  : in std_logic;

        poison_x  : out integer range 0 to GRID_WIDTH-1;
        poison_y  : out integer range 0 to GRID_HEIGHT-1;
        p1_poison : out std_logic;
        p2_poison : out std_logic
    );
end entity;

architecture rtl of poison_control is

    signal lfsr : std_logic_vector(9 downto 0) := SEED;

    signal poison_x_i : integer range 0 to GRID_WIDTH-1  := 10;
    signal poison_y_i : integer range 0 to GRID_HEIGHT-1 := 10;

    type state_t is (VISIBLE, HIDDEN);
    signal st : state_t := VISIBLE;

    signal hide_cnt : integer range 0 to HIDDEN_TICKS := 0;

    -- Border + random walls
    function is_wall_cell(
        x : integer;
        y : integer;
        w1_x0   : integer;
        w2_x0   : integer;
        w3_x0   : integer;
        w1_y0   : integer;
        w2_y0   : integer;
        w3_y0   : integer;
        w1_or   : std_logic;
        w2_or   : std_logic;
        w3_or   : std_logic;
        walls_s : std_logic
    ) return boolean is
    begin
        -- border
        if (x = 0) or (y = 0) or
           (x = GRID_WIDTH-1) or (y = GRID_HEIGHT-1) then
            return true;
        end if;

        -- solid random walls
        if walls_s = '1' then
            -- wall 1
            if w1_or = '0' then
                if (y = w1_y0) and (x >= w1_x0) and (x <= w1_x0 + 4) then
                    return true;
                end if;
            else
                if (x = w1_x0) and (y >= w1_y0) and (y <= w1_y0 + 4) then
                    return true;
                end if;
            end if;

            -- wall 2
            if w2_or = '0' then
                if (y = w2_y0) and (x >= w2_x0) and (x <= w2_x0 + 4) then
                    return true;
                end if;
            else
                if (x = w2_x0) and (y >= w2_y0) and (y <= w2_y0 + 4) then
                    return true;
                end if;
            end if;

            -- wall 3
            if w3_or = '0' then
                if (y = w3_y0) and (x >= w3_x0) and (x <= w3_x0 + 4) then
                    return true;
                end if;
            else
                if (x = w3_x0) and (y >= w3_y0) and (y <= w3_y0 + 4) then
                    return true;
                end if;
            end if;
        end if;

        return false;
    end function;

begin

    poison_x <= poison_x_i;
    poison_y <= poison_y_i;

    process(clk, rst)
        variable new_x    : integer range 0 to GRID_WIDTH-1;
        variable new_y    : integer range 0 to GRID_HEIGHT-1;
        variable x_raw    : integer;
        variable y_raw    : integer;
        variable nxt_lfsr : std_logic_vector(9 downto 0);
        variable p1_hit   : boolean;
        variable p2_hit   : boolean;
        variable j        : integer;
    begin
        if rst = '1' then
            lfsr        <= SEED;
            poison_x_i  <= 10;
            poison_y_i  <= 10;
            st          <= VISIBLE;
            hide_cnt    <= 0;
            p1_poison   <= '0';
            p2_poison   <= '0';
        elsif rising_edge(clk) then
            p1_poison <= '0';
            p2_poison <= '0';

            if game_tick = '1' then
                -- LFSR
                nxt_lfsr := lfsr(8 downto 0) & (lfsr(9) xor lfsr(6));
                lfsr     <= nxt_lfsr;

                case st is
                    when VISIBLE =>
                        p1_hit := (p1_head_x = poison_x_i) and (p1_head_y = poison_y_i);
                        p2_hit := (p2_head_x = poison_x_i) and (p2_head_y = poison_y_i);

                        if p1_hit or p2_hit then
                            if p1_hit then p1_poison <= '1'; end if;
                            if p2_hit then p2_poison <= '1'; end if;

                            -- new poison apple position: interior + avoid walls
                            x_raw := to_integer(unsigned(nxt_lfsr(5 downto 0)));
                            y_raw := to_integer(unsigned(nxt_lfsr(9 downto 6)));

                            new_x := 1 + (x_raw mod (GRID_WIDTH-2));
                            new_y := 1 + (y_raw mod (GRID_HEIGHT-2));

                            for j in 0 to 7 loop
                                exit when not is_wall_cell(
                                    new_x, new_y,
                                    w1_x0_i, w2_x0_i, w3_x0_i,
                                    w1_y0_i, w2_y0_i, w3_y0_i,
                                    w1_orient_i, w2_orient_i, w3_orient_i,
                                    walls_solid_i
                                );
                                new_x := 1 + ((new_x - 1 + 1) mod (GRID_WIDTH-2));
                                new_y := 1 + ((new_y - 1 + 1) mod (GRID_HEIGHT-2));
                            end loop;

                            poison_x_i <= new_x;
                            poison_y_i <= new_y;

                            st       <= HIDDEN;
                            hide_cnt <= 0;
                        end if;

                    when HIDDEN =>
                        if hide_cnt >= HIDDEN_TICKS then
                            st       <= VISIBLE;
                            hide_cnt <= 0;
                        else
                            hide_cnt <= hide_cnt + 1;
                        end if;
                end case;
            end if;
        end if;
    end process;

end architecture;
